////////////////////////////////////////////////////////////////////////////////////////////
module DATA_IN_VAR_RPI(
	//
	input [7:0] FPGA_TO_RPI_8BIT_01,
	input [7:0] FPGA_TO_RPI_8BIT_02,
	input [7:0] FPGA_TO_RPI_8BIT_03,
	input [7:0] FPGA_TO_RPI_8BIT_04,
	input [7:0] FPGA_TO_RPI_8BIT_05,
	input [7:0] FPGA_TO_RPI_8BIT_06,
	input [7:0] FPGA_TO_RPI_8BIT_07,
	input [7:0] FPGA_TO_RPI_8BIT_08,
	input [7:0] FPGA_TO_RPI_8BIT_09,
	//
	input [15:0] FPGA_TO_RPI_16BIT_01,
	input [15:0] FPGA_TO_RPI_16BIT_02,
	input [15:0] FPGA_TO_RPI_16BIT_03,
	input [15:0] FPGA_TO_RPI_16BIT_04,
	input [15:0] FPGA_TO_RPI_16BIT_05,
	input [15:0] FPGA_TO_RPI_16BIT_06,
	input [15:0] FPGA_TO_RPI_16BIT_07,
	input [15:0] FPGA_TO_RPI_16BIT_08,
	input [15:0] FPGA_TO_RPI_16BIT_09,
	input [15:0] FPGA_TO_RPI_16BIT_10,
	input [15:0] FPGA_TO_RPI_16BIT_11,
	input [15:0] FPGA_TO_RPI_16BIT_12,
	input [15:0] FPGA_TO_RPI_16BIT_13,
	input [15:0] FPGA_TO_RPI_16BIT_14,
	input [15:0] FPGA_TO_RPI_16BIT_15,
	input [15:0] FPGA_TO_RPI_16BIT_16,
	input [15:0] FPGA_TO_RPI_16BIT_17,
	input [15:0] FPGA_TO_RPI_16BIT_18,
	input [15:0] FPGA_TO_RPI_16BIT_19,
	input [15:0] FPGA_TO_RPI_16BIT_20,
	input [15:0] FPGA_TO_RPI_16BIT_21,
	input [15:0] FPGA_TO_RPI_16BIT_22,
	input [15:0] FPGA_TO_RPI_16BIT_23,
	input [15:0] FPGA_TO_RPI_16BIT_24,
	input [15:0] FPGA_TO_RPI_16BIT_25,
	input [15:0] FPGA_TO_RPI_16BIT_26,
	input [15:0] FPGA_TO_RPI_16BIT_27,
	//
	output [1023:0] DATA
	);
	//
	RPI_8BIT  rpi_8bit_01(FPGA_TO_RPI_8BIT_01[7:0],    DATA[015:008]);
	RPI_8BIT  rpi_8bit_02(FPGA_TO_RPI_8BIT_02[7:0],    DATA[023:016]);
	RPI_8BIT  rpi_8bit_03(FPGA_TO_RPI_8BIT_03[7:0],    DATA[031:024]);
	RPI_8BIT  rpi_8bit_04(FPGA_TO_RPI_8BIT_04[7:0],    DATA[039:032]);
	RPI_8BIT  rpi_8bit_05(FPGA_TO_RPI_8BIT_05[7:0],    DATA[047:040]);
	RPI_8BIT  rpi_8bit_06(FPGA_TO_RPI_8BIT_06[7:0],    DATA[055:048]);
	RPI_8BIT  rpi_8bit_07(FPGA_TO_RPI_8BIT_07[7:0],    DATA[063:056]);
	RPI_8BIT  rpi_8bit_08(FPGA_TO_RPI_8BIT_08[7:0],    DATA[071:064]);
	RPI_8BIT  rpi_8bit_09(FPGA_TO_RPI_8BIT_09[7:0],    DATA[079:072]);
	//
	RPI_16BIT rpi_16bit_01(FPGA_TO_RPI_16BIT_01[15:0], DATA[095:080]);
	RPI_16BIT rpi_16bit_02(FPGA_TO_RPI_16BIT_02[15:0], DATA[111:096]);
	RPI_16BIT rpi_16bit_03(FPGA_TO_RPI_16BIT_03[15:0], DATA[127:112]);
	RPI_16BIT rpi_16bit_04(FPGA_TO_RPI_16BIT_04[15:0], DATA[143:128]);
	RPI_16BIT rpi_16bit_05(FPGA_TO_RPI_16BIT_05[15:0], DATA[159:144]);
	RPI_16BIT rpi_16bit_06(FPGA_TO_RPI_16BIT_06[15:0], DATA[175:160]);
	RPI_16BIT rpi_16bit_07(FPGA_TO_RPI_16BIT_07[15:0], DATA[191:176]);
	RPI_16BIT rpi_16bit_08(FPGA_TO_RPI_16BIT_08[15:0], DATA[207:192]);
	RPI_16BIT rpi_16bit_09(FPGA_TO_RPI_16BIT_09[15:0], DATA[223:208]);
	RPI_16BIT rpi_16bit_10(FPGA_TO_RPI_16BIT_10[15:0], DATA[239:224]);
	RPI_16BIT rpi_16bit_11(FPGA_TO_RPI_16BIT_11[15:0], DATA[255:240]);
	RPI_16BIT rpi_16bit_12(FPGA_TO_RPI_16BIT_12[15:0], DATA[271:256]);
	RPI_16BIT rpi_16bit_13(FPGA_TO_RPI_16BIT_13[15:0], DATA[287:272]);
	RPI_16BIT rpi_16bit_14(FPGA_TO_RPI_16BIT_14[15:0], DATA[303:288]);
	RPI_16BIT rpi_16bit_15(FPGA_TO_RPI_16BIT_15[15:0], DATA[319:304]);
	RPI_16BIT rpi_16bit_16(FPGA_TO_RPI_16BIT_16[15:0], DATA[335:320]);
	RPI_16BIT rpi_16bit_17(FPGA_TO_RPI_16BIT_17[15:0], DATA[351:336]);
	RPI_16BIT rpi_16bit_18(FPGA_TO_RPI_16BIT_18[15:0], DATA[367:352]);
	RPI_16BIT rpi_16bit_19(FPGA_TO_RPI_16BIT_19[15:0], DATA[383:368]);
	RPI_16BIT rpi_16bit_20(FPGA_TO_RPI_16BIT_20[15:0], DATA[399:384]);
	RPI_16BIT rpi_16bit_21(FPGA_TO_RPI_16BIT_21[15:0], DATA[415:400]);
	RPI_16BIT rpi_16bit_22(FPGA_TO_RPI_16BIT_22[15:0], DATA[431:416]);
	RPI_16BIT rpi_16bit_23(FPGA_TO_RPI_16BIT_23[15:0], DATA[447:432]);
	RPI_16BIT rpi_16bit_24(FPGA_TO_RPI_16BIT_24[15:0], DATA[463:448]);
	RPI_16BIT rpi_16bit_25(FPGA_TO_RPI_16BIT_25[15:0], DATA[479:464]);
	RPI_16BIT rpi_16bit_26(FPGA_TO_RPI_16BIT_26[15:0], DATA[495:480]);
	RPI_16BIT rpi_16bit_27(FPGA_TO_RPI_16BIT_27[15:0], DATA[511:496]);
	//
endmodule
////////////////////////////////////////////////////////////////////////////////////////////
module DATA_OUT_VAR_RPI(
	//
	input [1023:0] DATA,
	//
	output [7:0] RPI_TO_FPGA_8BIT_01,
	output [7:0] RPI_TO_FPGA_8BIT_02,
	output [7:0] RPI_TO_FPGA_8BIT_03,
	output [7:0] RPI_TO_FPGA_8BIT_04,
	output [7:0] RPI_TO_FPGA_8BIT_05,
	output [7:0] RPI_TO_FPGA_8BIT_06,
	output [7:0] RPI_TO_FPGA_8BIT_07,
	output [7:0] RPI_TO_FPGA_8BIT_08,
	output [7:0] RPI_TO_FPGA_8BIT_09,
	output [7:0] RPI_TO_FPGA_8BIT_10,
	output [7:0] RPI_TO_FPGA_8BIT_11,
	output [7:0] RPI_TO_FPGA_8BIT_12,
	output [7:0] RPI_TO_FPGA_8BIT_13,
	output [7:0] RPI_TO_FPGA_8BIT_14,
	output [7:0] RPI_TO_FPGA_8BIT_15,
	output [7:0] RPI_TO_FPGA_8BIT_16,
	output [7:0] RPI_TO_FPGA_8BIT_17,
	output [7:0] RPI_TO_FPGA_8BIT_18,
	output [7:0] RPI_TO_FPGA_8BIT_19,
	output [7:0] RPI_TO_FPGA_8BIT_20,
	output [7:0] RPI_TO_FPGA_8BIT_21,
	output [7:0] RPI_TO_FPGA_8BIT_22,
	output [7:0] RPI_TO_FPGA_8BIT_23,
	output [7:0] RPI_TO_FPGA_8BIT_24,
	output [7:0] RPI_TO_FPGA_8BIT_25,
	output [7:0] RPI_TO_FPGA_8BIT_26,
	output [7:0] RPI_TO_FPGA_8BIT_27,
	output [7:0] RPI_TO_FPGA_8BIT_28,
	output [7:0] RPI_TO_FPGA_8BIT_29,
	output [7:0] RPI_TO_FPGA_8BIT_30,
	output [7:0] RPI_TO_FPGA_8BIT_31,
	output [7:0] RPI_TO_FPGA_8BIT_32,
	output [7:0] RPI_TO_FPGA_8BIT_33,
	//
	output [15:0] RPI_TO_FPGA_16BIT_01,
	output [15:0] RPI_TO_FPGA_16BIT_02,
	output [15:0] RPI_TO_FPGA_16BIT_03,
	output [15:0] RPI_TO_FPGA_16BIT_04,
	output [15:0] RPI_TO_FPGA_16BIT_05,
	output [15:0] RPI_TO_FPGA_16BIT_06,
	output [15:0] RPI_TO_FPGA_16BIT_07,
	output [15:0] RPI_TO_FPGA_16BIT_08,
	output [15:0] RPI_TO_FPGA_16BIT_09,
	output [15:0] RPI_TO_FPGA_16BIT_10,
	output [15:0] RPI_TO_FPGA_16BIT_11,
	output [15:0] RPI_TO_FPGA_16BIT_12,
	output [15:0] RPI_TO_FPGA_16BIT_13,
	output [15:0] RPI_TO_FPGA_16BIT_14,
	output [15:0] RPI_TO_FPGA_16BIT_15,
	output [15:0] RPI_TO_FPGA_16BIT_16,
	output [15:0] RPI_TO_FPGA_16BIT_17,
	output [15:0] RPI_TO_FPGA_16BIT_18,
	output [15:0] RPI_TO_FPGA_16BIT_19,
	output [15:0] RPI_TO_FPGA_16BIT_20,
	output [15:0] RPI_TO_FPGA_16BIT_21,
	output [15:0] RPI_TO_FPGA_16BIT_22,
	output [15:0] RPI_TO_FPGA_16BIT_23,
	output [15:0] RPI_TO_FPGA_16BIT_24,
	output [15:0] RPI_TO_FPGA_16BIT_25,
	output [15:0] RPI_TO_FPGA_16BIT_26,
	output [15:0] RPI_TO_FPGA_16BIT_27
	);
	//
	RPI_8BIT rpi_8bit_01(DATA[015:008],   RPI_TO_FPGA_8BIT_01[7:0]);
	RPI_8BIT rpi_8bit_02(DATA[023:016],   RPI_TO_FPGA_8BIT_02[7:0]);
	RPI_8BIT rpi_8bit_03(DATA[031:024],   RPI_TO_FPGA_8BIT_03[7:0]);
	RPI_8BIT rpi_8bit_04(DATA[039:032],   RPI_TO_FPGA_8BIT_04[7:0]);
	RPI_8BIT rpi_8bit_05(DATA[047:040],   RPI_TO_FPGA_8BIT_05[7:0]);
	RPI_8BIT rpi_8bit_06(DATA[055:048],   RPI_TO_FPGA_8BIT_06[7:0]);
	RPI_8BIT rpi_8bit_07(DATA[063:056],   RPI_TO_FPGA_8BIT_07[7:0]);
	RPI_8BIT rpi_8bit_08(DATA[071:064],   RPI_TO_FPGA_8BIT_08[7:0]);
	RPI_8BIT rpi_8bit_09(DATA[079:072],   RPI_TO_FPGA_8BIT_09[7:0]);
	RPI_8BIT rpi_8bit_10(DATA[087:080],   RPI_TO_FPGA_8BIT_10[7:0]);
	RPI_8BIT rpi_8bit_11(DATA[095:088],   RPI_TO_FPGA_8BIT_11[7:0]);
	RPI_8BIT rpi_8bit_12(DATA[103:096],   RPI_TO_FPGA_8BIT_12[7:0]);
	RPI_8BIT rpi_8bit_13(DATA[111:104],   RPI_TO_FPGA_8BIT_13[7:0]);
	RPI_8BIT rpi_8bit_14(DATA[119:112],   RPI_TO_FPGA_8BIT_14[7:0]);
	RPI_8BIT rpi_8bit_15(DATA[127:120],   RPI_TO_FPGA_8BIT_15[7:0]);
	RPI_8BIT rpi_8bit_16(DATA[135:128],   RPI_TO_FPGA_8BIT_16[7:0]);
	RPI_8BIT rpi_8bit_17(DATA[143:136],   RPI_TO_FPGA_8BIT_17[7:0]);
	RPI_8BIT rpi_8bit_18(DATA[151:144],   RPI_TO_FPGA_8BIT_18[7:0]);
	RPI_8BIT rpi_8bit_19(DATA[159:152],   RPI_TO_FPGA_8BIT_19[7:0]);
	RPI_8BIT rpi_8bit_20(DATA[167:160],   RPI_TO_FPGA_8BIT_20[7:0]);
	RPI_8BIT rpi_8bit_21(DATA[175:168],   RPI_TO_FPGA_8BIT_21[7:0]);
	RPI_8BIT rpi_8bit_22(DATA[183:176],   RPI_TO_FPGA_8BIT_22[7:0]);
	RPI_8BIT rpi_8bit_23(DATA[191:184],   RPI_TO_FPGA_8BIT_23[7:0]);
	RPI_8BIT rpi_8bit_24(DATA[199:192],   RPI_TO_FPGA_8BIT_24[7:0]);
	RPI_8BIT rpi_8bit_25(DATA[207:200],   RPI_TO_FPGA_8BIT_25[7:0]);
	RPI_8BIT rpi_8bit_26(DATA[215:208],   RPI_TO_FPGA_8BIT_26[7:0]);
	RPI_8BIT rpi_8bit_27(DATA[223:216],   RPI_TO_FPGA_8BIT_27[7:0]);
	RPI_8BIT rpi_8bit_28(DATA[231:224],   RPI_TO_FPGA_8BIT_28[7:0]);
	RPI_8BIT rpi_8bit_29(DATA[239:232],   RPI_TO_FPGA_8BIT_29[7:0]);
	RPI_8BIT rpi_8bit_30(DATA[247:240],   RPI_TO_FPGA_8BIT_30[7:0]);
	RPI_8BIT rpi_8bit_31(DATA[255:248],   RPI_TO_FPGA_8BIT_31[7:0]);
	RPI_8BIT rpi_8bit_32(DATA[263:256],   RPI_TO_FPGA_8BIT_32[7:0]);
	RPI_8BIT rpi_8bit_33(DATA[271:264],   RPI_TO_FPGA_8BIT_33[7:0]);
	//
	RPI_16BIT rpi_16bit_01(DATA[287:272], RPI_TO_FPGA_16BIT_01[15:0]);
	RPI_16BIT rpi_16bit_02(DATA[303:288], RPI_TO_FPGA_16BIT_02[15:0]);
	RPI_16BIT rpi_16bit_03(DATA[319:304], RPI_TO_FPGA_16BIT_03[15:0]);
	RPI_16BIT rpi_16bit_04(DATA[335:320], RPI_TO_FPGA_16BIT_04[15:0]);
	RPI_16BIT rpi_16bit_05(DATA[351:336], RPI_TO_FPGA_16BIT_05[15:0]);
	RPI_16BIT rpi_16bit_06(DATA[367:352], RPI_TO_FPGA_16BIT_06[15:0]);
	RPI_16BIT rpi_16bit_07(DATA[383:368], RPI_TO_FPGA_16BIT_07[15:0]);
	RPI_16BIT rpi_16bit_08(DATA[399:384], RPI_TO_FPGA_16BIT_08[15:0]);
	RPI_16BIT rpi_16bit_09(DATA[415:400], RPI_TO_FPGA_16BIT_09[15:0]);
	RPI_16BIT rpi_16bit_10(DATA[431:416], RPI_TO_FPGA_16BIT_10[15:0]);
	RPI_16BIT rpi_16bit_11(DATA[447:432], RPI_TO_FPGA_16BIT_11[15:0]);
	RPI_16BIT rpi_16bit_12(DATA[463:448], RPI_TO_FPGA_16BIT_12[15:0]);
	RPI_16BIT rpi_16bit_13(DATA[479:464], RPI_TO_FPGA_16BIT_13[15:0]);
	RPI_16BIT rpi_16bit_14(DATA[495:480], RPI_TO_FPGA_16BIT_14[15:0]);
	RPI_16BIT rpi_16bit_15(DATA[511:496], RPI_TO_FPGA_16BIT_15[15:0]);
	RPI_16BIT rpi_16bit_16(DATA[527:512], RPI_TO_FPGA_16BIT_16[15:0]);
	RPI_16BIT rpi_16bit_17(DATA[543:528], RPI_TO_FPGA_16BIT_17[15:0]);
	RPI_16BIT rpi_16bit_18(DATA[559:544], RPI_TO_FPGA_16BIT_18[15:0]);
	RPI_16BIT rpi_16bit_19(DATA[575:560], RPI_TO_FPGA_16BIT_19[15:0]);
	RPI_16BIT rpi_16bit_20(DATA[591:576], RPI_TO_FPGA_16BIT_20[15:0]);
	RPI_16BIT rpi_16bit_21(DATA[607:592], RPI_TO_FPGA_16BIT_21[15:0]);
	RPI_16BIT rpi_16bit_22(DATA[623:608], RPI_TO_FPGA_16BIT_22[15:0]);
	RPI_16BIT rpi_16bit_23(DATA[639:624], RPI_TO_FPGA_16BIT_23[15:0]);
	RPI_16BIT rpi_16bit_24(DATA[655:640], RPI_TO_FPGA_16BIT_24[15:0]);
	RPI_16BIT rpi_16bit_25(DATA[671:656], RPI_TO_FPGA_16BIT_25[15:0]);
	RPI_16BIT rpi_16bit_26(DATA[687:672], RPI_TO_FPGA_16BIT_26[15:0]);
	RPI_16BIT rpi_16bit_27(DATA[703:688], RPI_TO_FPGA_16BIT_27[15:0]);
	//
	//Prozessabbild: 88 Bytes
endmodule
////////////////////////////////////////////////////////////////////////////////////////////
module RPI_32BIT(
	input [31:0] IN,
	output [31:0] OUT
	);
	//
	RPI_8BIT rpi_8bit_1(IN[31:24], OUT[31:24]);
	RPI_8BIT rpi_8bit_2(IN[23:16], OUT[23:16]);
	RPI_8BIT rpi_8bit_3(IN[15:08], OUT[15:08]);
	RPI_8BIT rpi_8bit_4(IN[07:00], OUT[07:00]);
	//
endmodule
//
module RPI_16BIT(
	input [15:0] IN,
	output [15:0] OUT
	);
	//
	RPI_8BIT rpi_8bit_1(IN[15:08], OUT[15:08]);
	RPI_8BIT rpi_8bit_2(IN[07:00], OUT[07:00]);
	
	//
endmodule
//
module RPI_8BIT(
	input [7:0] IN,
	output [7:0] OUT
	);
	//	
	assign OUT[0] = IN[7];	
	assign OUT[1] = IN[6];	
	assign OUT[2] = IN[5];	
	assign OUT[3] = IN[4];	
	assign OUT[4] = IN[3];	
	assign OUT[5] = IN[2];	
	assign OUT[6] = IN[1];
	assign OUT[7] = IN[0];
	//
endmodule
////////////////////////////////////////////////////////////////////////////////////////////
