
module ISSP (
	source);	

	output	[0:0]	source;
endmodule
