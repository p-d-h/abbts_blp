module CONST_8 (
	output [7:0] OUT
	);
	//	
	parameter VALUE = 8'd1;
	//
	assign OUT = VALUE;
endmodule